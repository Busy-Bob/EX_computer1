library verilog;
use verilog.vl_types.all;
entity test_computer_vlg_vec_tst is
end test_computer_vlg_vec_tst;
